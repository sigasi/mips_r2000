library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity ROM_atpgHamming is
	port( clk,rst : in std_logic;
			do_ROM  : out std_logic_vector(37 downto 0));
end ROM_atpgHamming;

architecture Behavioral of ROM_atpgHamming is

begin


end Behavioral;

