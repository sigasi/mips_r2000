library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use ieee.std_logic_unsigned.all;

entity ROM_mem_vectors is
	port( clk,rst : in std_logic;
			do : out std_logic_vector(63 downto 0));
end ROM_mem_vectors;

architecture Behavioral of ROM_mem_vectors is

type ROM is array (0 to 87) of std_logic_vector(63 downto 0);
signal mem : Rom := ("0100001000001110001001001000000000000000000001100000000000000100",           --ATPG VECTORS FOR TESTING
							"0100110110110101001001001001000010111001010111000000000000000111",
                     "0111110101000100000001001110000010001111010100101000011000001000",
							"0010010110110000001001000001000011010001111011000000000010110010",	
							"1000001000110101000001000001000010000000000000000000011000000000",
							"0101000001000110001001001111011010010001111000000000000000000100",
							"0100000001001000110101110111011011101000000000000000000000000000",
							"1100000000000001001001111111111000000000000000000000011011011000",
							"0110001100111000111001000011010011011010011010101001110111101000",
							"0101001000101001000001001000000000010000000000000000010000100100",
							"0101010000001110101001001001000010011010000000000000000011000000",
							"0100001000000010010011010110010100000001111100000100010000100100",
							"0000000101011011010001000101000001001000000000101100011111100001",
							"0111100001000110001000000001000001110010000000000000000110000010",
							"1010000111110101001001001000000011010001111000000000000000100000",
							"1010001101001100001110000001000000001101001101010000000000110010",
							"1100000001000001001000001111001100000000000000000000000001100100",
							"0000010010001010010010000000100000111001101001111100110110110001",
							"0000001000110101001001001001001011100000000000000000001100000000",
							"0101001001001001001001111111010100000110010010001000000001111001",
							"0001100110100001000001110001000010111011101000000011000000001000",
							"0001001000000000000001000001110111000000000000000000000000000001",
							"0000110001000001001000000010010100000000100000000011100000000000",
							"0001100111000111000101000101000011010011010101001110000010000101",
							"1111010100001000000001001000100000111101000110101100000000000100",
							"1001111000001001000101000000000000011100000000000001001011001000",
							"0100001000001110001001001001000100000000000000110000000000000100",
							"0101000000001001001110101001000000101010000000000110000000000000",
							"1110000001111100001011001011111110000000100011001011001111100110",
							"1010000110011100011100100001001000111101001101010100111010110010",
							"0001011101110001001001001110000001010110010000100000110000000010",
							"0100100101000101101100110100000100000011000000011100100111010110",
							"0100110101010111010100001001000000111110111110010011000010110010",
							"1011101001001000001001001000000010010000000000000000000000000011",
							"1000001000000001000110101000000011000000000011000000000000000000",
							"1111001001000001000001110010111100000000000011110001101111001001",
							"0100001001001000000000000110000100110000000000000000000000000100",
							"0010001100001000001000000110000010001010000011000000000000001000",
							"0111101001000000000000001000110011010011100000000000000000000100",
							"0101001001000000000101000001100100000000000001010100111110010010",
							"1111001001001001001001110011011000000000100000000111010000111111",
							"1000100101100101000101000001000010111111111010000000000010000101",
							"1000001111100001011000000000000001111111000100110100000000000100",
							"0100110001001000001001000110011000000000000000000001101001100000",
							"0000001000001001110100110111111000011000000000000000000000000100",
							"0101001000110000001001110110010100000000001101000000000001111111",
							"1110000010011101010010000011111110001010111100100111100001001001",
							"0000100111000010110000100111110001010101100011111101001010100101",
							"0100110001000001000110010010111000100000000011100000000001111111",
							"0010001111100001001001000101000000100100011001011000001000010010",
							"1001001110000001000001001000000001000000000000000000000001100100",
							"0001001000110100110010010011010100111000000000000000000101110100",
							"0010101010001111001000001000001000110010110100000000000000001100",
							"1001001000001001001000110101001011000000000110000000000000000000",
							"1100001000101001001001001001000011111011110000000000000000000111",
							"1011000100111010100001001000001010111101111001001100000010110010",
							"1001000111110000101100110001000010010010001100101100111000111010",
							"1110001111001110011010110110111001000001110100100000100100011001",
							"1001111101000100010110010011111100100111110110101111111011001111",
							"0100001001111011110110011111110101000000000000111000111000110010",
							"0001001011011000110100100001000001101000111101101001000000000001",
							"0100000000001001000110101000000010000000000110000000000000000000",
							"0100000001001000010111111111001100000100000000000000100100000111",
							"0101000001001110000010111111111101100100000000000000000001111101",
							"0100101001000001000000000110001010000000000000000000000010110100",
							"0101001000000001001001001000110001110000000000000000000000010000",
							"0000110011010001001000110001001001011101110110100000000110000010",
							"0101001001001001001001001001000100000000000000000000000000010101",
							"0001000000110001001001110010010110010001111000000000000000000100",
							"0001010001101001100000000000100011100001101001101000010000000000",
							"0100000110000001111110011111011100100001101100000000011100110111",
							"0111000001000001110001000000000010000010000000000000110000000010",
							"1000010100011010011100001000000010111000011010011010100000000100",
							"0000101100001000000001001001110000010001111110000000000000000010",
							"1111001000110001001001001001001000101100000000000000000000001001",
							"0000000111000000001000001111010000000000000001111000000000000100",
							"0011111101010001000000011110100111100011110101001010000000001110",
							"0100001000001110000001001001100000000000000110000000000000000000",
							"0100000110001111111000101101110010000000000000000011001101101000",
							"1001000000000001110101000000000010000000000000001100000000000000",
							"1100001011011000001110000000000001110011000011000000000011001000",
							"0110101000000001000000000001000100000000000000000001100000001000",
							"0100001001001001000001110001000100000001100000000000000000000001",
							"1001000001000110001000001001000001000000000000000011000000000001",
							"0000101001000000000000001000001010000000000000000000000000001000",
							"0011010010011000101000001110100011000010101100101000011000000000",
							"1001101001001100011101010110001011100001010110010100110001110001",
							"0100001000001000110000001000100000000000110000000000000000000100");
						
signal addr : std_logic_vector(6 downto 0) := "0000000";

begin
	process(clk)
	begin
		if(rising_edge(clk))then
			do <= mem( to_integer(unsigned(addr)));
			
--			if(rst = '1') then
--				addr <= "0000";
--			else
--				addr <= addr + "0001";
--			end if;
		end if;
	end process;
	process(clk)
	begin
		if(rising_edge(clk))then
			if(rst = '1') then
				addr <= "0000000";
			else
				addr <= addr + "0000001";
			end if;
		end if;
	
	end process;
	

end Behavioral;